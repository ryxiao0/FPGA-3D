module z_buffer(
    input wire clk_in,
    input wire rst_in,
    output logic [23:0] pixel_color
);

    

endmodule