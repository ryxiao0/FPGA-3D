module scaling
    (
        input wire clk_in,
        input wire rst_in,
        output logic valid_out
    );

    logic x;

endmodule