$date
   Thu Dec  7 12:10:04 2023
$end
$version
  2023.1
$end
$timescale
  1ps
$end
$scope module tri_proj_tb $end
$var reg 1 ! clk $end
$var reg 1 " rst $end
$var reg 32 # x_in [31:0] $end
$var reg 32 $ y_in [31:0] $end
$var reg 32 % z_in [31:0] $end
$var reg 1 & v_in $end
$var reg 9 ' x [8:0] $end
$var reg 9 ( y [8:0] $end
$var reg 9 ) z [8:0] $end
$var reg 1 * v_out $end
$scope module uut $end
$var wire 1 + clk_in $end
$var wire 1 , rst_in $end
$var wire 1 - obj_done_in $end
$var wire 1 . valid_in $end
$var reg 9 ' x [8:0] $end
$var reg 9 ( y [8:0] $end
$var reg 9 ) z [8:0] $end
$var reg 1 * valid_out $end
$var reg 1 / obj_done_out $end
$var reg 32 0 state $end
$var reg 32 1 rec_in [31:0] $end
$var reg 32 2 rec_out [31:0] $end
$var reg 1 3 rec_v_in $end
$var reg 1 4 rec_v_out $end
$var reg 32 5 mult_a_in [31:0] $end
$var reg 32 6 mult_b_in [31:0] $end
$var reg 32 7 mult_out [31:0] $end
$var reg 1 8 mult_v_in $end
$var reg 1 9 mult_v_out $end
$var reg 32 : round_in [31:0] $end
$var reg 16 ; round_out [15:0] $end
$var reg 1 < round_v_in $end
$var reg 1 = round_v_out $end
$var reg 32 > x_f [31:0] $end
$var reg 32 ? y_f [31:0] $end
$var reg 32 @ z_f [31:0] $end
$var reg 10 A shift [9:0] $end
$scope module rec $end
$var wire 1 + aclk $end
$var wire 1 B s_axis_a_tvalid $end
$var wire 1 C s_axis_a_tready $end
$var wire 32 D s_axis_a_tdata [31:0] $end
$var wire 1 E m_axis_result_tvalid $end
$var wire 1 F m_axis_result_tready $end
$var wire 32 G m_axis_result_tdata [31:0] $end
$upscope $end
$scope module pro $end
$var wire 1 + aclk $end
$var wire 1 H s_axis_a_tvalid $end
$var wire 1 I s_axis_a_tready $end
$var wire 32 J s_axis_a_tdata [31:0] $end
$var wire 1 K s_axis_b_tvalid $end
$var wire 1 L s_axis_b_tready $end
$var wire 32 M s_axis_b_tdata [31:0] $end
$var wire 1 N m_axis_result_tvalid $end
$var wire 1 O m_axis_result_tready $end
$var wire 32 P m_axis_result_tdata [31:0] $end
$upscope $end
$scope module round $end
$var wire 1 + aclk $end
$var wire 1 Q s_axis_a_tvalid $end
$var wire 1 R s_axis_a_tready $end
$var wire 32 S s_axis_a_tdata [31:0] $end
$var wire 1 T m_axis_result_tvalid $end
$var wire 1 U m_axis_result_tready $end
$var wire 16 V m_axis_result_tdata [15:0] $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
0!
0"
bx #
bx $
bx %
x&
bx '
bx (
bx )
x*
0+
0,
z-
x.
z/
b0 0
bx 1
b0 2
x3
04
bx 5
bx 6
b0 7
x8
09
bx :
b0 ;
x<
0=
bx >
bx ?
bx @
b10110100 A
xB
1C
bx D
0E
1F
b0 G
xH
1I
bx J
xK
1L
bx M
0N
1O
b0 P
xQ
1R
bx S
0T
1U
b0 V
$end
#5000
1!
1"
0*
1+
1,
b1111110100000000000000000000000 2
b1111110100000000000000000000000 G
#10000
0!
0+
#15000
1!
0"
1+
0,
#20000
0!
0+
#25000
1!
b1000000110000000000000000000000 #
b1000000110000000000000000000000 $
b1000000110000000000000000000000 %
1&
1+
1.
b1 0
b1000000110000000000000000000000 5
b111110010011001100110011001101 6
b1000000000000000000000000000000 7
18
b1000000110000000000000000000000 @
1H
b1000000110000000000000000000000 J
1K
b111110010011001100110011001101 M
b1000000000000000000000000000000 P
#30000
0!
0+
#35000
1!
0&
1+
0.
08
0H
0K
#40000
0!
0+
#45000
1!
1+
b100000000000000 ;
b110110100 A
b100000000000000 V
#50000
0!
0+
#55000
1!
1+
b0 ;
b10110100 A
b0 V
#60000
0!
0+
#65000
1!
1+
b0 7
b0 P
#70000
0!
0+
#75000
1!
1+
#80000
0!
0+
#85000
1!
1+
#90000
0!
0+
#95000
1!
1+
#100000
0!
0+
#105000
1!
1+
#110000
0!
0+
#115000
1!
1+
b111111100110011001100110011010 7
19
1N
b111111100110011001100110011010 P
#120000
0!
0+
#125000
1!
1+
b10 0
b111111100110011001100110011010 1
13
09
1B
b111111100110011001100110011010 D
0N
#130000
0!
0+
#135000
1!
1+
03
0B
#140000
0!
0+
#145000
1!
1+
#150000
0!
0+
#155000
1!
1+
#160000
0!
0+
#165000
1!
1+
#170000
0!
0+
#175000
1!
1+
#180000
0!
0+
#185000
1!
1+
#190000
0!
0+
#195000
1!
1+
#200000
0!
0+
#205000
1!
1+
#210000
0!
0+
#215000
1!
1+
#220000
0!
0+
#225000
1!
1+
#230000
0!
0+
#235000
1!
1+
#240000
0!
0+
#245000
1!
1+
#250000
0!
0+
#255000
1!
1+
#260000
0!
0+
#265000
1!
1+
#270000
0!
0+
#275000
1!
1+
#280000
0!
0+
#285000
1!
1+
b1111111100000000000000000000000 2
b1111111100000000000000000000000 G
#290000
0!
0+
#295000
1!
1+
#300000
0!
0+
#305000
1!
1+
#310000
0!
0+
#315000
1!
1+
#320000
0!
0+
#325000
1!
1+
#330000
0!
0+
#335000
1!
1+
#340000
0!
0+
#345000
1!
1+
#350000
0!
0+
#355000
1!
1+
#360000
0!
0+
#365000
1!
1+
#370000
0!
0+
#375000
1!
1+
#380000
0!
0+
#385000
1!
1+
#390000
0!
0+
#395000
1!
1+
#400000
0!
0+
#405000
1!
1+
#410000
0!
0+
#415000
1!
1+
#420000
0!
0+
#425000
1!
1+
b111111010101010101010101010101 2
14
1E
b111111010101010101010101010101 G
#430000
0!
0+
#435000
1!
1+
b11 0
04
b111111010101010101010101010101 5
b1000000110000000000000000000000 6
18
0E
1H
b111111010101010101010101010101 J
1K
b1000000110000000000000000000000 M
#440000
0!
0+
#445000
1!
1+
08
0H
0K
#450000
0!
0+
#455000
1!
1+
#460000
0!
0+
#465000
1!
1+
#470000
0!
0+
#475000
1!
1+
#480000
0!
0+
#485000
1!
1+
#490000
0!
0+
#495000
1!
1+
#500000
0!
0+
#505000
1!
1+
#510000
0!
0+
#515000
1!
1+
#520000
0!
0+
#525000
1!
1+
b1000000101000000000000000000000 7
19
1N
b1000000101000000000000000000000 P
#530000
0!
0+
#535000
1!
1+
b100 0
18
09
b1000000101000000000000000000000 >
1H
1K
0N
#540000
0!
0+
#545000
1!
1+
08
0H
0K
#550000
0!
0+
#555000
1!
1+
#560000
0!
0+
#565000
1!
1+
#570000
0!
0+
#575000
1!
1+
#580000
0!
0+
#585000
1!
1+
#590000
0!
0+
#595000
1!
1+
#600000
0!
0+
#605000
1!
1+
#610000
0!
0+
#615000
1!
1+
#620000
0!
0+
#625000
1!
1+
19
1N
#630000
0!
0+
#635000
1!
1+
b101 0
b1000011001101000000000000000000 5
b1000000101000000000000000000000 6
18
09
b1000000101000000000000000000000 ?
1H
b1000011001101000000000000000000 J
1K
b1000000101000000000000000000000 M
0N
#640000
0!
0+
#645000
1!
1+
08
0H
0K
#650000
0!
0+
#655000
1!
1+
#660000
0!
0+
#665000
1!
1+
#670000
0!
0+
#675000
1!
1+
#680000
0!
0+
#685000
1!
1+
#690000
0!
0+
#695000
1!
1+
#700000
0!
0+
#705000
1!
1+
#710000
0!
0+
#715000
1!
1+
#720000
0!
0+
#725000
1!
1+
b1000100011000010000000000000000 7
19
1N
b1000100011000010000000000000000 P
#730000
0!
0+
#735000
1!
1+
b110 0
09
b1000100011000010000000000000000 :
1<
0N
1Q
b1000100011000010000000000000000 S
#740000
0!
0+
#745000
1!
1+
0<
0Q
#750000
0!
0+
#755000
1!
1+
#760000
0!
0+
#765000
1!
1+
#770000
0!
0+
#775000
1!
1+
#780000
0!
0+
#785000
1!
1+
#790000
0!
0+
#795000
1!
1+
#800000
0!
0+
#805000
1!
1+
b111111111111111 ;
1=
b1010110011 A
1T
b111111111111111 V
#810000
0!
0+
#815000
1!
b10110011 '
1+
b111 0
18
0=
1H
1K
0T
#820000
0!
0+
#825000
1!
1+
08
0H
0K
#830000
0!
0+
#835000
1!
1+
#840000
0!
0+
#845000
1!
1+
#850000
0!
0+
#855000
1!
1+
#860000
0!
0+
#865000
1!
1+
#870000
0!
0+
#875000
1!
1+
#880000
0!
0+
#885000
1!
1+
#890000
0!
0+
#895000
1!
1+
#900000
0!
0+
#905000
1!
1+
19
1N
#910000
0!
0+
#915000
1!
1+
b1000 0
09
1<
0N
1Q
#920000
0!
0+
#925000
1!
1+
0<
0Q
#930000
0!
0+
#935000
1!
1+
#940000
0!
0+
#945000
1!
1+
#950000
0!
0+
#955000
1!
1+
#960000
0!
0+
#965000
1!
1+
#970000
0!
0+
#975000
1!
1+
#980000
0!
0+
#985000
1!
1+
1=
1T
#990000
0!
0+
#995000
1!
b10110011 (
1+
b1001 0
b1000000110000000000000000000000 6
18
0=
1H
1K
b1000000110000000000000000000000 M
0T
#1000000
0!
0+
