$date
   Wed Dec  6 23:49:11 2023
$end
$version
  2023.1
$end
$timescale
  1ps
$end
$scope module tri_proj_tb $end
$var reg 1 ! clk $end
$var reg 1 " rst $end
$var reg 32 # x_in [31:0] $end
$var reg 32 $ y_in [31:0] $end
$var reg 32 % z_in [31:0] $end
$var reg 1 & v_in $end
$var reg 32 ' x [31:0] $end
$var reg 32 ( y [31:0] $end
$var reg 1 ) v_out $end
$scope module uut $end
$var wire 1 * clk_in $end
$var wire 1 + rst_in $end
$var wire 1 , valid_in $end
$var reg 1 ) valid_out $end
$var reg 32 - state $end
$var reg 32 . rec_in [31:0] $end
$var reg 32 / rec_out [31:0] $end
$var reg 1 0 rec_v_in $end
$var reg 1 1 rec_v_out $end
$var reg 32 2 mult_a_in [31:0] $end
$var reg 32 3 mult_b_in [31:0] $end
$var reg 32 4 mult_out [31:0] $end
$var reg 1 5 mult_v_in $end
$var reg 1 6 mult_v_out $end
$scope module rec $end
$var wire 1 * aclk $end
$var wire 1 7 s_axis_a_tvalid $end
$var wire 1 8 s_axis_a_tready $end
$var wire 32 9 s_axis_a_tdata [31:0] $end
$var wire 1 : m_axis_result_tvalid $end
$var wire 1 ; m_axis_result_tready $end
$var wire 32 < m_axis_result_tdata [31:0] $end
$upscope $end
$scope module pro $end
$var wire 1 * aclk $end
$var wire 1 = s_axis_a_tvalid $end
$var wire 1 > s_axis_a_tready $end
$var wire 32 ? s_axis_a_tdata [31:0] $end
$var wire 1 @ s_axis_b_tvalid $end
$var wire 1 A s_axis_b_tready $end
$var wire 32 B s_axis_b_tdata [31:0] $end
$var wire 1 C m_axis_result_tvalid $end
$var wire 1 D m_axis_result_tready $end
$var wire 32 E m_axis_result_tdata [31:0] $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
0!
0"
bx #
bx $
bx %
x&
bx '
bx (
x)
0*
0+
x,
b0 -
bx .
b0 /
x0
01
bx 2
bx 3
b0 4
x5
06
x7
18
bx 9
0:
1;
b0 <
x=
1>
bx ?
x@
1A
bx B
0C
1D
b0 E
$end
#5000
1!
1"
0)
1*
1+
b1111110100000000000000000000000 /
b1111110100000000000000000000000 <
#10000
0!
0*
#15000
1!
0"
1*
0+
#20000
0!
0*
#25000
1!
b1000000110000000000000000000000 #
b1000000110000000000000000000000 $
b1000000110000000000000000000000 %
1&
1*
1,
b1 -
b1000000110000000000000000000000 2
b111110010011001100110011001101 3
b1000000000000000000000000000000 4
15
1=
b1000000110000000000000000000000 ?
1@
b111110010011001100110011001101 B
b1000000000000000000000000000000 E
#30000
0!
0*
#35000
1!
0&
1*
0,
05
0=
0@
#40000
0!
0*
#45000
1!
1*
#50000
0!
0*
#55000
1!
1*
#60000
0!
0*
#65000
1!
1*
b0 4
b0 E
#70000
0!
0*
#75000
1!
1*
#80000
0!
0*
#85000
1!
1*
#90000
0!
0*
#95000
1!
1*
#100000
0!
0*
#105000
1!
1*
#110000
0!
0*
#115000
1!
1*
b111111100110011001100110011010 4
16
1C
b111111100110011001100110011010 E
#120000
0!
0*
#125000
1!
1*
b10 -
b111111100110011001100110011010 .
10
06
17
b111111100110011001100110011010 9
0C
#130000
0!
0*
#135000
1!
1*
00
07
#140000
0!
0*
#145000
1!
1*
#150000
0!
0*
#155000
1!
1*
#160000
0!
0*
#165000
1!
1*
#170000
0!
0*
#175000
1!
1*
#180000
0!
0*
#185000
1!
1*
#190000
0!
0*
#195000
1!
1*
#200000
0!
0*
#205000
1!
1*
#210000
0!
0*
#215000
1!
1*
#220000
0!
0*
#225000
1!
1*
#230000
0!
0*
#235000
1!
1*
#240000
0!
0*
#245000
1!
1*
#250000
0!
0*
#255000
1!
1*
#260000
0!
0*
#265000
1!
1*
#270000
0!
0*
#275000
1!
1*
#280000
0!
0*
#285000
1!
1*
b1111111100000000000000000000000 /
b1111111100000000000000000000000 <
#290000
0!
0*
#295000
1!
1*
#300000
0!
0*
#305000
1!
1*
#310000
0!
0*
#315000
1!
1*
#320000
0!
0*
#325000
1!
1*
#330000
0!
0*
#335000
1!
1*
#340000
0!
0*
#345000
1!
1*
#350000
0!
0*
#355000
1!
1*
#360000
0!
0*
#365000
1!
1*
#370000
0!
0*
#375000
1!
1*
#380000
0!
0*
#385000
1!
1*
#390000
0!
0*
#395000
1!
1*
#400000
0!
0*
#405000
1!
1*
#410000
0!
0*
#415000
1!
1*
#420000
0!
0*
#425000
1!
1*
b111111010101010101010101010101 /
11
1:
b111111010101010101010101010101 <
#430000
0!
0*
#435000
1!
1*
b11 -
01
b111111010101010101010101010101 2
b1000000110000000000000000000000 3
15
0:
1=
b111111010101010101010101010101 ?
1@
b1000000110000000000000000000000 B
#440000
0!
0*
#445000
1!
1*
05
0=
0@
#450000
0!
0*
#455000
1!
1*
#460000
0!
0*
#465000
1!
1*
#470000
0!
0*
#475000
1!
1*
#480000
0!
0*
#485000
1!
1*
#490000
0!
0*
#495000
1!
1*
#500000
0!
0*
#505000
1!
1*
#510000
0!
0*
#515000
1!
1*
#520000
0!
0*
#525000
1!
1*
b1000000101000000000000000000000 4
16
1C
b1000000101000000000000000000000 E
#530000
0!
0*
#535000
1!
b1000000101000000000000000000000 '
1*
b100 -
15
06
1=
1@
0C
#540000
0!
0*
#545000
1!
1*
05
0=
0@
#550000
0!
0*
#555000
1!
1*
#560000
0!
0*
#565000
1!
1*
#570000
0!
0*
#575000
1!
1*
#580000
0!
0*
#585000
1!
1*
#590000
0!
0*
#595000
1!
1*
#600000
0!
0*
#605000
1!
1*
#610000
0!
0*
#615000
1!
1*
#620000
0!
0*
#625000
1!
1*
16
1C
#630000
0!
0*
#635000
1!
b1000000101000000000000000000000 (
1)
1*
b0 -
06
0C
#640000
0!
0*
#645000
1!
0)
1*
#650000
0!
0*
#655000
1!
1*
#660000
0!
0*
#665000
1!
1*
#670000
0!
0*
#675000
1!
1*
#680000
0!
0*
#685000
1!
1*
#690000
0!
0*
#695000
1!
1*
#700000
0!
0*
#705000
1!
1*
#710000
0!
0*
#715000
1!
1*
#720000
0!
0*
#725000
1!
1*
#730000
0!
0*
#735000
1!
1*
#740000
0!
0*
#745000
1!
1*
#750000
0!
0*
#755000
1!
1*
#760000
0!
0*
#765000
1!
1*
#770000
0!
0*
#775000
1!
1*
#780000
0!
0*
#785000
1!
1*
#790000
0!
0*
#795000
1!
1*
#800000
0!
0*
#805000
1!
1*
#810000
0!
0*
#815000
1!
1*
#820000
0!
0*
#825000
1!
1*
#830000
0!
0*
#835000
1!
1*
#840000
0!
0*
#845000
1!
1*
#850000
0!
0*
#855000
1!
1*
#860000
0!
0*
#865000
1!
1*
#870000
0!
0*
#875000
1!
1*
#880000
0!
0*
#885000
1!
1*
#890000
0!
0*
#895000
1!
1*
#900000
0!
0*
#905000
1!
1*
#910000
0!
0*
#915000
1!
1*
#920000
0!
0*
#925000
1!
1*
#930000
0!
0*
#935000
1!
1*
#940000
0!
0*
#945000
1!
1*
#950000
0!
0*
#955000
1!
1*
#960000
0!
0*
#965000
1!
1*
#970000
0!
0*
#975000
1!
1*
#980000
0!
0*
#985000
1!
1*
#990000
0!
0*
#995000
1!
1*
#1000000
0!
0*
