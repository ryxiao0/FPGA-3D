$date
   Wed Dec 13 21:57:22 2023
$end
$version
  2023.1
$end
$timescale
  1ps
$end
$scope module transformation_tb $end
$var reg 1 ! clk $end
$var reg 1 " rst $end
$var reg 32 # x_in [31:0] $end
$var reg 32 $ y_in [31:0] $end
$var reg 32 % z_in [31:0] $end
$var reg 1 & v_in $end
$var reg 32 ' x [31:0] $end
$var reg 32 ( y [31:0] $end
$var reg 32 ) z [31:0] $end
$var reg 32 * w [31:0] $end
$var reg 1 + v_out $end
$var reg 32 , distance [31:0] $end
$var reg 1 - ready_out $end
$var reg 1 . ready_in $end
$var reg 1 / obj_done_in $end
$var reg 1 0 obj_done_out $end
$scope module uut $end
$var wire 1 1 clk_in $end
$var wire 1 2 rst_in $end
$var wire 32 3 distance [31:0] $end
$var wire 32 4 scale [31:0] $end
$var wire 5 5 pitch [4:0] $end
$var wire 5 6 roll [4:0] $end
$var wire 5 7 yaw [4:0] $end
$var wire 1 8 obj_done_in $end
$var wire 1 9 valid_in $end
$var reg 1 + valid_out $end
$var reg 1 0 obj_done_out $end
$var reg 1 - ready_out $end
$var wire 1 : ready_in $end
$var reg 32 ; state $end
$var reg 32 < add_a_in [31:0] $end
$var reg 32 = add_b_in [31:0] $end
$var reg 32 > add_out [31:0] $end
$var reg 1 ? add_v_in $end
$var reg 1 @ add_v_out $end
$var reg 32 A mult_a_in [31:0] $end
$var reg 32 B mult_b_in [31:0] $end
$var reg 32 C mult_out [31:0] $end
$var reg 1 D mult_v_in $end
$var reg 1 E mult_v_out $end
$scope module add $end
$var wire 1 1 aclk $end
$var wire 1 F s_axis_a_tvalid $end
$var wire 1 G s_axis_a_tready $end
$var wire 32 H s_axis_a_tdata [31:0] $end
$var wire 1 I s_axis_b_tvalid $end
$var wire 1 J s_axis_b_tready $end
$var wire 32 K s_axis_b_tdata [31:0] $end
$var wire 1 L m_axis_result_tvalid $end
$var wire 1 M m_axis_result_tready $end
$var wire 32 N m_axis_result_tdata [31:0] $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
0!
0"
bx #
bx $
bx %
x&
bx '
bx (
bx )
bx *
x+
bx ,
x-
x.
x/
x0
01
02
bx 3
bz 4
bz 5
bz 6
bz 7
x8
x9
x:
b0 ;
bx <
bx =
bx >
x?
0@
bx A
bx B
bx C
xD
xE
xF
1G
bx H
xI
1J
bx K
0L
1M
bx N
$end
#5000
1!
1"
0+
11
12
b0 >
b0 N
#10000
0!
01
#15000
1!
0"
11
02
#20000
0!
b111111100000000000000000000000 #
b111111100000000000000000000000 $
b111111100000000000000000000000 %
1&
b1000001001000000000000000000000 ,
1.
1/
10
01
b1000001001000000000000000000000 3
18
19
1:
#25000
1!
11
b1 ;
b111111100000000000000000000000 <
b1000001001000000000000000000000 =
1?
1F
b111111100000000000000000000000 H
1I
b1000001001000000000000000000000 K
#30000
0!
0&
01
09
#35000
1!
11
0?
0F
0I
#40000
0!
01
#45000
1!
11
#50000
0!
01
#55000
1!
11
#60000
0!
01
#65000
1!
11
#70000
0!
01
#75000
1!
11
#80000
0!
01
#85000
1!
11
#90000
0!
01
#95000
1!
11
b100000000000000000000000 >
b100000000000000000000000 N
#100000
0!
01
#105000
1!
11
b0 >
b0 N
#110000
0!
01
#115000
1!
11
#120000
0!
01
#125000
1!
11
#130000
0!
01
#135000
1!
11
#140000
0!
01
#145000
1!
11
b1000001001100000000000000000000 >
1@
1L
b1000001001100000000000000000000 N
#150000
0!
01
#155000
1!
b111111100000000000000000000000 '
b111111100000000000000000000000 (
b1000001001100000000000000000000 )
b111111100000000000000000000000 *
1+
11
b0 ;
0@
0L
#160000
0!
01
#165000
1!
0+
11
#170000
0!
01
#175000
1!
11
#180000
0!
01
#185000
1!
11
#190000
0!
01
#195000
1!
11
#200000
0!
01
#205000
1!
11
#210000
0!
01
#215000
1!
11
#220000
0!
01
#225000
1!
11
#230000
0!
01
#235000
1!
11
#240000
0!
01
#245000
1!
11
#250000
0!
01
#255000
1!
11
#260000
0!
01
#265000
1!
11
#270000
0!
01
#275000
1!
11
#280000
0!
01
#285000
1!
11
#290000
0!
01
#295000
1!
11
#300000
0!
01
#305000
1!
11
#310000
0!
01
#315000
1!
11
#320000
0!
01
#325000
1!
11
#330000
0!
01
#335000
1!
11
#340000
0!
01
#345000
1!
11
#350000
0!
01
#355000
1!
11
#360000
0!
01
#365000
1!
11
#370000
0!
01
#375000
1!
11
#380000
0!
01
#385000
1!
11
#390000
0!
01
#395000
1!
11
#400000
0!
01
#405000
1!
11
#410000
0!
01
#415000
1!
11
#420000
0!
01
#425000
1!
11
#430000
0!
01
#435000
1!
11
#440000
0!
01
#445000
1!
11
#450000
0!
01
#455000
1!
11
#460000
0!
01
#465000
1!
11
#470000
0!
01
#475000
1!
11
#480000
0!
01
#485000
1!
11
#490000
0!
01
#495000
1!
11
#500000
0!
01
#505000
1!
11
#510000
0!
01
#515000
1!
11
#520000
0!
01
#525000
1!
11
#530000
0!
01
#535000
1!
11
#540000
0!
01
#545000
1!
11
#550000
0!
01
#555000
1!
11
#560000
0!
01
#565000
1!
11
#570000
0!
01
#575000
1!
11
#580000
0!
01
#585000
1!
11
#590000
0!
01
#595000
1!
11
#600000
0!
01
#605000
1!
11
#610000
0!
01
#615000
1!
11
#620000
0!
01
#625000
1!
11
#630000
0!
01
#635000
1!
11
#640000
0!
01
#645000
1!
11
#650000
0!
01
#655000
1!
11
#660000
0!
01
#665000
1!
11
#670000
0!
01
#675000
1!
11
#680000
0!
01
#685000
1!
11
#690000
0!
01
#695000
1!
11
#700000
0!
01
#705000
1!
11
#710000
0!
01
#715000
1!
11
#720000
0!
01
#725000
1!
11
#730000
0!
01
#735000
1!
11
#740000
0!
01
#745000
1!
11
#750000
0!
01
#755000
1!
11
#760000
0!
01
#765000
1!
11
#770000
0!
01
#775000
1!
11
#780000
0!
01
#785000
1!
11
#790000
0!
01
#795000
1!
11
#800000
0!
01
#805000
1!
11
#810000
0!
01
#815000
1!
11
#820000
0!
01
#825000
1!
11
#830000
0!
01
#835000
1!
11
#840000
0!
01
#845000
1!
11
#850000
0!
01
#855000
1!
11
#860000
0!
01
#865000
1!
11
#870000
0!
01
#875000
1!
11
#880000
0!
01
#885000
1!
11
#890000
0!
01
#895000
1!
11
#900000
0!
01
#905000
1!
11
#910000
0!
01
#915000
1!
11
#920000
0!
01
#925000
1!
11
#930000
0!
01
#935000
1!
11
#940000
0!
01
#945000
1!
11
#950000
0!
01
#955000
1!
11
#960000
0!
01
#965000
1!
11
#970000
0!
01
#975000
1!
11
#980000
0!
01
#985000
1!
11
#990000
0!
01
#995000
1!
11
#1000000
0!
01
