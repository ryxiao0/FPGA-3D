module rotation
    (
        input wire clk_in,
        input wire rst_in,
        input wire [31:0] pitch,
        input wire [31:0] roll,
        input wire [31:0] yaw,
        input wire [31:0] vertex [4:0]
    );

    logic x;

endmodule