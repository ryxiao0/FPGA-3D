module rasterizer (
    input wire clk_in,
    input wire rst_in,
    output logic triangle [2:0]
);



endmodule