$date
   Wed Dec  6 13:40:09 2023
$end
$version
  2023.1
$end
$timescale
  1ps
$end
$scope module transformation_tb $end
$var reg 1 ! clk $end
$var reg 1 " rst $end
$var reg 1 # v_in $end
$var reg 32 $ x [31:0] $end
$var reg 32 % y [31:0] $end
$var reg 32 & z [31:0] $end
$var reg 32 ' w [31:0] $end
$var reg 1 ( v_out $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
0!
0"
x#
bx $
bx %
bx &
bx '
x(
$end
#5000
1!
1"
#10000
0!
#15000
1!
0"
#20000
0!
1#
#25000
1!
#30000
0!
0#
#35000
1!
#40000
0!
#45000
1!
#50000
0!
#55000
1!
#60000
0!
#65000
1!
#70000
0!
#75000
1!
#80000
0!
#85000
1!
#90000
0!
#95000
1!
#100000
0!
#105000
1!
#110000
0!
#115000
1!
#120000
0!
#125000
1!
#130000
0!
#135000
1!
#140000
0!
#145000
1!
#150000
0!
#155000
1!
#160000
0!
#165000
1!
#170000
0!
#175000
1!
#180000
0!
#185000
1!
#190000
0!
#195000
1!
#200000
0!
#205000
1!
#210000
0!
#215000
1!
#220000
0!
#225000
1!
#230000
0!
#235000
1!
#240000
0!
#245000
1!
#250000
0!
#255000
1!
#260000
0!
#265000
1!
#270000
0!
#275000
1!
#280000
0!
#285000
1!
#290000
0!
#295000
1!
#300000
0!
#305000
1!
#310000
0!
#315000
1!
#320000
0!
#325000
1!
#330000
0!
#335000
1!
#340000
0!
#345000
1!
#350000
0!
#355000
1!
#360000
0!
#365000
1!
#370000
0!
#375000
1!
#380000
0!
#385000
1!
#390000
0!
#395000
1!
#400000
0!
#405000
1!
#410000
0!
#415000
1!
#420000
0!
#425000
1!
#430000
0!
#435000
1!
#440000
0!
#445000
1!
#450000
0!
#455000
1!
#460000
0!
#465000
1!
#470000
0!
#475000
1!
#480000
0!
#485000
1!
#490000
0!
#495000
1!
#500000
0!
#505000
1!
#510000
0!
#515000
1!
#520000
0!
#525000
1!
#530000
0!
#535000
1!
#540000
0!
#545000
1!
#550000
0!
#555000
1!
#560000
0!
#565000
1!
#570000
0!
#575000
1!
#580000
0!
#585000
1!
#590000
0!
#595000
1!
#600000
0!
#605000
1!
#610000
0!
#615000
1!
#620000
0!
#625000
1!
#630000
0!
#635000
1!
#640000
0!
#645000
1!
#650000
0!
#655000
1!
#660000
0!
#665000
1!
#670000
0!
#675000
1!
#680000
0!
#685000
1!
#690000
0!
#695000
1!
#700000
0!
#705000
1!
#710000
0!
#715000
1!
#720000
0!
#725000
1!
#730000
0!
#735000
1!
#740000
0!
#745000
1!
#750000
0!
#755000
1!
#760000
0!
#765000
1!
#770000
0!
#775000
1!
#780000
0!
#785000
1!
#790000
0!
#795000
1!
#800000
0!
#805000
1!
#810000
0!
#815000
1!
#820000
0!
#825000
1!
#830000
0!
#835000
1!
#840000
0!
#845000
1!
#850000
0!
#855000
1!
#860000
0!
#865000
1!
#870000
0!
#875000
1!
#880000
0!
#885000
1!
#890000
0!
#895000
1!
#900000
0!
#905000
1!
#910000
0!
#915000
1!
#920000
0!
#925000
1!
#930000
0!
#935000
1!
#940000
0!
#945000
1!
#950000
0!
#955000
1!
#960000
0!
#965000
1!
#970000
0!
#975000
1!
#980000
0!
#985000
1!
#990000
0!
#995000
1!
#1000000
0!
