$date
   Wed Dec  6 13:55:45 2023
$end
$version
  2023.1
$end
$timescale
  1ps
$end
$scope module transformation_tb $end
$var reg 1 ! clk $end
$var reg 1 " rst $end
$var reg 32 # x_in [31:0] $end
$var reg 32 $ y_in [31:0] $end
$var reg 32 % z_in [31:0] $end
$var reg 1 & v_in $end
$var reg 32 ' x [31:0] $end
$var reg 32 ( y [31:0] $end
$var reg 32 ) z [31:0] $end
$var reg 32 * w [31:0] $end
$var reg 1 + v_out $end
$scope module uut $end
$var wire 1 , clk_in $end
$var wire 1 - rst_in $end
$var wire 2 . sel [1:0] $end
$var wire 32 / scale [31:0] $end
$var wire 5 0 pitch [4:0] $end
$var wire 5 1 roll [4:0] $end
$var wire 5 2 yaw [4:0] $end
$var wire 1 3 valid_in $end
$var reg 1 + valid_out $end
$var reg 32 4 state $end
$var reg 32 5 add_a_in [31:0] $end
$var reg 32 6 add_b_in [31:0] $end
$var reg 32 7 add_out [31:0] $end
$var reg 1 8 add_v_in $end
$var reg 1 9 add_v_out $end
$var reg 32 : mult_a_in [31:0] $end
$var reg 32 ; mult_b_in [31:0] $end
$var reg 32 < mult_out [31:0] $end
$var reg 1 = mult_v_in $end
$var reg 1 > mult_v_out $end
$scope module add $end
$var wire 1 , aclk $end
$var wire 1 ? s_axis_a_tvalid $end
$var wire 1 @ s_axis_a_tready $end
$var wire 32 A s_axis_a_tdata [31:0] $end
$var wire 1 B s_axis_b_tvalid $end
$var wire 1 C s_axis_b_tready $end
$var wire 32 D s_axis_b_tdata [31:0] $end
$var wire 1 E m_axis_result_tvalid $end
$var wire 1 F m_axis_result_tready $end
$var wire 32 G m_axis_result_tdata [31:0] $end
$upscope $end
$scope module mult $end
$var wire 1 , aclk $end
$var wire 1 H s_axis_a_tvalid $end
$var wire 1 I s_axis_a_tready $end
$var wire 32 J s_axis_a_tdata [31:0] $end
$var wire 1 K s_axis_b_tvalid $end
$var wire 1 L s_axis_b_tready $end
$var wire 32 M s_axis_b_tdata [31:0] $end
$var wire 1 N m_axis_result_tvalid $end
$var wire 1 O m_axis_result_tready $end
$var wire 32 P m_axis_result_tdata [31:0] $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
0!
0"
bx #
bx $
bx %
x&
bx '
bx (
bx )
bx *
x+
0,
0-
bz .
bz /
bz 0
bz 1
bz 2
x3
b0 4
bx 5
bx 6
bx 7
x8
09
bx :
bx ;
b0 <
x=
0>
x?
1@
bx A
xB
1C
bx D
0E
1F
bx G
xH
1I
bx J
xK
1L
bx M
0N
1O
b0 P
$end
#5000
1!
1"
0+
1,
1-
b0 7
b0 G
#10000
0!
0,
#15000
1!
0"
1,
0-
#20000
0!
1&
b0 '
b0 (
b0 )
0,
13
#25000
1!
1,
b1 4
b1010 6
18
b1000000000000000000000000000000 <
1?
1B
b1010 D
b1000000000000000000000000000000 P
#30000
0!
0&
0,
03
#35000
1!
1,
08
0?
0B
#40000
0!
0,
#45000
1!
1,
#50000
0!
0,
#55000
1!
1,
#60000
0!
0,
#65000
1!
1,
b0 <
b0 P
#70000
0!
0,
#75000
1!
1,
#80000
0!
0,
#85000
1!
1,
#90000
0!
0,
#95000
1!
1,
b100000000000000000000000 7
b100000000000000000000000 G
#100000
0!
0,
#105000
1!
1,
b0 7
b0 G
#110000
0!
0,
#115000
1!
1,
#120000
0!
0,
#125000
1!
1,
#130000
0!
0,
#135000
1!
1,
#140000
0!
0,
#145000
1!
1,
19
1E
#150000
0!
0,
#155000
1!
b111111100000000000000000000000 *
1+
1,
b0 4
09
0E
#160000
0!
0,
#165000
1!
0+
1,
#170000
0!
0,
#175000
1!
1,
#180000
0!
0,
#185000
1!
1,
#190000
0!
0,
#195000
1!
1,
#200000
0!
0,
#205000
1!
1,
#210000
0!
0,
#215000
1!
1,
#220000
0!
0,
#225000
1!
1,
#230000
0!
0,
#235000
1!
1,
#240000
0!
0,
#245000
1!
1,
#250000
0!
0,
#255000
1!
1,
#260000
0!
0,
#265000
1!
1,
#270000
0!
0,
#275000
1!
1,
#280000
0!
0,
#285000
1!
1,
#290000
0!
0,
#295000
1!
1,
#300000
0!
0,
#305000
1!
1,
#310000
0!
0,
#315000
1!
1,
#320000
0!
0,
#325000
1!
1,
#330000
0!
0,
#335000
1!
1,
#340000
0!
0,
#345000
1!
1,
#350000
0!
0,
#355000
1!
1,
#360000
0!
0,
#365000
1!
1,
#370000
0!
0,
#375000
1!
1,
#380000
0!
0,
#385000
1!
1,
#390000
0!
0,
#395000
1!
1,
#400000
0!
0,
#405000
1!
1,
#410000
0!
0,
#415000
1!
1,
#420000
0!
0,
#425000
1!
1,
#430000
0!
0,
#435000
1!
1,
#440000
0!
0,
#445000
1!
1,
#450000
0!
0,
#455000
1!
1,
#460000
0!
0,
#465000
1!
1,
#470000
0!
0,
#475000
1!
1,
#480000
0!
0,
#485000
1!
1,
#490000
0!
0,
#495000
1!
1,
#500000
0!
0,
#505000
1!
1,
#510000
0!
0,
#515000
1!
1,
#520000
0!
0,
#525000
1!
1,
#530000
0!
0,
#535000
1!
1,
#540000
0!
0,
#545000
1!
1,
#550000
0!
0,
#555000
1!
1,
#560000
0!
0,
#565000
1!
1,
#570000
0!
0,
#575000
1!
1,
#580000
0!
0,
#585000
1!
1,
#590000
0!
0,
#595000
1!
1,
#600000
0!
0,
#605000
1!
1,
#610000
0!
0,
#615000
1!
1,
#620000
0!
0,
#625000
1!
1,
#630000
0!
0,
#635000
1!
1,
#640000
0!
0,
#645000
1!
1,
#650000
0!
0,
#655000
1!
1,
#660000
0!
0,
#665000
1!
1,
#670000
0!
0,
#675000
1!
1,
#680000
0!
0,
#685000
1!
1,
#690000
0!
0,
#695000
1!
1,
#700000
0!
0,
#705000
1!
1,
#710000
0!
0,
#715000
1!
1,
#720000
0!
0,
#725000
1!
1,
#730000
0!
0,
#735000
1!
1,
#740000
0!
0,
#745000
1!
1,
#750000
0!
0,
#755000
1!
1,
#760000
0!
0,
#765000
1!
1,
#770000
0!
0,
#775000
1!
1,
#780000
0!
0,
#785000
1!
1,
#790000
0!
0,
#795000
1!
1,
#800000
0!
0,
#805000
1!
1,
#810000
0!
0,
#815000
1!
1,
#820000
0!
0,
#825000
1!
1,
#830000
0!
0,
#835000
1!
1,
#840000
0!
0,
#845000
1!
1,
#850000
0!
0,
#855000
1!
1,
#860000
0!
0,
#865000
1!
1,
#870000
0!
0,
#875000
1!
1,
#880000
0!
0,
#885000
1!
1,
#890000
0!
0,
#895000
1!
1,
#900000
0!
0,
#905000
1!
1,
#910000
0!
0,
#915000
1!
1,
#920000
0!
0,
#925000
1!
1,
#930000
0!
0,
#935000
1!
1,
#940000
0!
0,
#945000
1!
1,
#950000
0!
0,
#955000
1!
1,
#960000
0!
0,
#965000
1!
1,
#970000
0!
0,
#975000
1!
1,
#980000
0!
0,
#985000
1!
1,
#990000
0!
0,
#995000
1!
1,
#1000000
0!
0,
